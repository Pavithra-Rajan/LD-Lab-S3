
module not_gate(I,O);
	input I;
	output O;
	nand(O,I,I);
endmodule
